library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package aes_tboxes_pkg is
  subtype u8  is std_logic_vector(7 downto 0);
  subtype u32 is std_logic_vector(31 downto 0);

  type tbox32_t is array (0 to 255) of u32;
  type tbox8_t  is array (0 to 255) of u8;

  -- Encryption T-boxes (from OpenSSL Te0..Te3)
  constant Te0 : tbox32_t;
  constant Te1 : tbox32_t;
  constant Te2 : tbox32_t;
  constant Te3 : tbox32_t;
  -- S-box for final round (equivalent to Te4)
  constant Te4 : tbox8_t;

  -- Decryption T-boxes (Td0..Td3) and Td4 (inverse S)
  constant Td0 : tbox32_t;
  constant Td1 : tbox32_t;
  constant Td2 : tbox32_t;
  constant Td3 : tbox32_t;
  constant Td4 : tbox8_t;

end package;

package body aes_tboxes_pkg is

  -- OpenSSL AES T-boxes
  constant Te0 : tbox32_t := (
    x"c66363a5", x"f87c7c84", x"ee777799", x"f67b7b8d",
    x"fff2f20d", x"d66b6bbd", x"de6f6fb1", x"91c5c554",
    x"60303050", x"02010103", x"ce6767a9", x"562b2b7d",
    x"e7fefe19", x"b5d7d762", x"4dababe6", x"ec76769a",
    x"8fcaca45", x"1f82829d", x"89c9c940", x"fa7d7d87",
    x"effafa15", x"b25959eb", x"8e4747c9", x"fbf0f00b",
    x"41adadec", x"b3d4d467", x"5fa2a2fd", x"45afafea",
    x"239c9cbf", x"53a4a4f7", x"e4727296", x"9bc0c05b",
    x"75b7b7c2", x"e1fdfd1c", x"3d9393ae", x"4c26266a",
    x"6c36365a", x"7e3f3f41", x"f5f7f702", x"83cccc4f",
    x"6834345c", x"51a5a5f4", x"d1e5e534", x"f9f1f108",
    x"e2717193", x"abd8d873", x"62313153", x"2a15153f",
    x"0804040c", x"95c7c752", x"46232365", x"9dc3c35e",
    x"30181828", x"379696a1", x"0a05050f", x"2f9a9ab5",
    x"0e070709", x"24121236", x"1b80809b", x"dfe2e23d",
    x"cdebeb26", x"4e272769", x"7fb2b2cd", x"ea75759f",
    x"1209091b", x"1d83839e", x"582c2c74", x"341a1a2e",
    x"361b1b2d", x"dc6e6eb2", x"b45a5aee", x"5ba0a0fb",
    x"a45252f6", x"763b3b4d", x"b7d6d661", x"7db3b3ce",
    x"5229297b", x"dde3e33e", x"5e2f2f71", x"13848497",
    x"a65353f5", x"b9d1d168", x"00000000", x"c1eded2c",
    x"40202060", x"e3fcfc1f", x"79b1b1c8", x"b65b5bed",
    x"d46a6abe", x"8dcbcb46", x"67bebed9", x"7239394b",
    x"944a4ade", x"984c4cd4", x"b05858e8", x"85cfcf4a",
    x"bbd0d06b", x"c5efef2a", x"4faaaae5", x"edfbfb16",
    x"864343c5", x"9a4d4dd7", x"66333355", x"11858594",
    x"8a4545cf", x"e9f9f910", x"04020206", x"fe7f7f81",
    x"a05050f0", x"783c3c44", x"259f9fba", x"4ba8a8e3",
    x"a25151f3", x"5da3a3fe", x"804040c0", x"058f8f8a",
    x"3f9292ad", x"219d9dbc", x"70383848", x"f1f5f504",
    x"63bcbcdf", x"77b6b6c1", x"afdada75", x"42212163",
    x"20101030", x"e5ffff1a", x"fdf3f30e", x"bfd2d26d",
    x"81cdcd4c", x"180c0c14", x"26131335", x"c3ecec2f",
    x"be5f5fe1", x"359797a2", x"884444cc", x"2e171739",
    x"93c4c457", x"55a7a7f2", x"fc7e7e82", x"7a3d3d47",
    x"c86464ac", x"ba5d5de7", x"3219192b", x"e6737395",
    x"c06060a0", x"19818198", x"9e4f4fd1", x"a3dcdc7f",
    x"44222266", x"542a2a7e", x"3b9090ab", x"0b888883",
    x"8c4646ca", x"c7eeee29", x"6bb8b8d3", x"2814143c",
    x"a7dede79", x"bc5e5ee2", x"160b0b1d", x"addbdb76",
    x"dbe0e03b", x"64323256", x"743a3a4e", x"140a0a1e",
    x"924949db", x"0c06060a", x"4824246c", x"b85c5ce4",
    x"9fc2c25d", x"bdd3d36e", x"43acacef", x"c46262a6",
    x"399191a8", x"319595a4", x"d3e4e437", x"f279798b",
    x"d5e7e732", x"8bc8c843", x"6e373759", x"da6d6db7",
    x"018d8d8c", x"b1d5d564", x"9c4e4ed2", x"49a9a9e0",
    x"d86c6cb4", x"ac5656fa", x"f3f4f407", x"cfeaea25",
    x"ca6565af", x"f47a7a8e", x"47aeaee9", x"10080818",
    x"6fbabad5", x"f0787888", x"4a25256f", x"5c2e2e72",
    x"381c1c24", x"57a6a6f1", x"73b4b4c7", x"97c6c651",
    x"cbe8e823", x"a1dddd7c", x"e874749c", x"3e1f1f21",
    x"964b4bdd", x"61bdbddc", x"0d8b8b86", x"0f8a8a85",
    x"e0707090", x"7c3e3e42", x"71b5b5c4", x"cc6666aa",
    x"904848d8", x"06030305", x"f7f6f601", x"1c0e0e12",
    x"c26161a3", x"6a35355f", x"ae5757f9", x"69b9b9d0",
    x"17868691", x"99c1c158", x"3a1d1d27", x"279e9eb9",
    x"d9e1e138", x"ebf8f813", x"2b9898b3", x"22111133",
    x"d26969bb", x"a9d9d970", x"078e8e89", x"339494a7",
    x"2d9b9bb6", x"3c1e1e22", x"15878792", x"c9e9e920",
    x"87cece49", x"aa5555ff", x"50282878", x"a5dfdf7a",
    x"038c8c8f", x"59a1a1f8", x"09898980", x"1a0d0d17",
    x"65bfbfda", x"d7e6e631", x"844242c6", x"d06868b8",
    x"824141c3", x"299999b0", x"5a2d2d77", x"1e0f0f11",
    x"7bb0b0cb", x"a85454fc", x"6dbbbbd6", x"2c16163a"
  );
  constant Te1 : tbox32_t := (
    x"a5c66363", x"84f87c7c", x"99ee7777", x"8df67b7b",
    x"0dfff2f2", x"bdd66b6b", x"b1de6f6f", x"5491c5c5",
    x"50603030", x"03020101", x"a9ce6767", x"7d562b2b",
    x"19e7fefe", x"62b5d7d7", x"e64dabab", x"9aec7676",
    x"458fcaca", x"9d1f8282", x"4089c9c9", x"87fa7d7d",
    x"15effafa", x"ebb25959", x"c98e4747", x"0bfbf0f0",
    x"ec41adad", x"67b3d4d4", x"fd5fa2a2", x"ea45afaf",
    x"bf239c9c", x"f753a4a4", x"96e47272", x"5b9bc0c0",
    x"c275b7b7", x"1ce1fdfd", x"ae3d9393", x"6a4c2626",
    x"5a6c3636", x"417e3f3f", x"02f5f7f7", x"4f83cccc",
    x"5c683434", x"f451a5a5", x"34d1e5e5", x"08f9f1f1",
    x"93e27171", x"73abd8d8", x"53623131", x"3f2a1515",
    x"0c080404", x"5295c7c7", x"65462323", x"5e9dc3c3",
    x"28301818", x"a1379696", x"0f0a0505", x"b52f9a9a",
    x"090e0707", x"36241212", x"9b1b8080", x"3ddfe2e2",
    x"26cdebeb", x"694e2727", x"cd7fb2b2", x"9fea7575",
    x"1b120909", x"9e1d8383", x"74582c2c", x"2e341a1a",
    x"2d361b1b", x"b2dc6e6e", x"eeb45a5a", x"fb5ba0a0",
    x"f6a45252", x"4d763b3b", x"61b7d6d6", x"ce7db3b3",
    x"7b522929", x"3edde3e3", x"715e2f2f", x"97138484",
    x"f5a65353", x"68b9d1d1", x"00000000", x"2cc1eded",
    x"60402020", x"1fe3fcfc", x"c879b1b1", x"edb65b5b",
    x"bed46a6a", x"468dcbcb", x"d967bebe", x"4b723939",
    x"de944a4a", x"d4984c4c", x"e8b05858", x"4a85cfcf",
    x"6bbbd0d0", x"2ac5efef", x"e54faaaa", x"16edfbfb",
    x"c5864343", x"d79a4d4d", x"55663333", x"94118585",
    x"cf8a4545", x"10e9f9f9", x"06040202", x"81fe7f7f",
    x"f0a05050", x"44783c3c", x"ba259f9f", x"e34ba8a8",
    x"f3a25151", x"fe5da3a3", x"c0804040", x"8a058f8f",
    x"ad3f9292", x"bc219d9d", x"48703838", x"04f1f5f5",
    x"df63bcbc", x"c177b6b6", x"75afdada", x"63422121",
    x"30201010", x"1ae5ffff", x"0efdf3f3", x"6dbfd2d2",
    x"4c81cdcd", x"14180c0c", x"35261313", x"2fc3ecec",
    x"e1be5f5f", x"a2359797", x"cc884444", x"392e1717",
    x"5793c4c4", x"f255a7a7", x"82fc7e7e", x"477a3d3d",
    x"acc86464", x"e7ba5d5d", x"2b321919", x"95e67373",
    x"a0c06060", x"98198181", x"d19e4f4f", x"7fa3dcdc",
    x"66442222", x"7e542a2a", x"ab3b9090", x"830b8888",
    x"ca8c4646", x"29c7eeee", x"d36bb8b8", x"3c281414",
    x"79a7dede", x"e2bc5e5e", x"1d160b0b", x"76addbdb",
    x"3bdbe0e0", x"56643232", x"4e743a3a", x"1e140a0a",
    x"db924949", x"0a0c0606", x"6c482424", x"e4b85c5c",
    x"5d9fc2c2", x"6ebdd3d3", x"ef43acac", x"a6c46262",
    x"a8399191", x"a4319595", x"37d3e4e4", x"8bf27979",
    x"32d5e7e7", x"438bc8c8", x"596e3737", x"b7da6d6d",
    x"8c018d8d", x"64b1d5d5", x"d29c4e4e", x"e049a9a9",
    x"b4d86c6c", x"faac5656", x"07f3f4f4", x"25cfeaea",
    x"afca6565", x"8ef47a7a", x"e947aeae", x"18100808",
    x"d56fbaba", x"88f07878", x"6f4a2525", x"725c2e2e",
    x"24381c1c", x"f157a6a6", x"c773b4b4", x"5197c6c6",
    x"23cbe8e8", x"7ca1dddd", x"9ce87474", x"213e1f1f",
    x"dd964b4b", x"dc61bdbd", x"860d8b8b", x"850f8a8a",
    x"90e07070", x"427c3e3e", x"c471b5b5", x"aacc6666",
    x"d8904848", x"05060303", x"01f7f6f6", x"121c0e0e",
    x"a3c26161", x"5f6a3535", x"f9ae5757", x"d069b9b9",
    x"91178686", x"5899c1c1", x"273a1d1d", x"b9279e9e",
    x"38d9e1e1", x"13ebf8f8", x"b32b9898", x"33221111",
    x"bbd26969", x"70a9d9d9", x"89078e8e", x"a7339494",
    x"b62d9b9b", x"223c1e1e", x"92158787", x"20c9e9e9",
    x"4987cece", x"ffaa5555", x"78502828", x"7aa5dfdf",
    x"8f038c8c", x"f859a1a1", x"80098989", x"171a0d0d",
    x"da65bfbf", x"31d7e6e6", x"c6844242", x"b8d06868",
    x"c3824141", x"b0299999", x"775a2d2d", x"111e0f0f",
    x"cb7bb0b0", x"fca85454", x"d66dbbbb", x"3a2c1616"
  );
  constant Te2 : tbox32_t := (
    x"63a5c663", x"7c84f87c", x"7799ee77", x"7b8df67b",
    x"f20dfff2", x"6bbdd66b", x"6fb1de6f", x"c55491c5",
    x"30506030", x"01030201", x"67a9ce67", x"2b7d562b",
    x"fe19e7fe", x"d762b5d7", x"abe64dab", x"769aec76",
    x"ca458fca", x"829d1f82", x"c94089c9", x"7d87fa7d",
    x"fa15effa", x"59ebb259", x"47c98e47", x"f00bfbf0",
    x"adec41ad", x"d467b3d4", x"a2fd5fa2", x"afea45af",
    x"9cbf239c", x"a4f753a4", x"7296e472", x"c05b9bc0",
    x"b7c275b7", x"fd1ce1fd", x"93ae3d93", x"266a4c26",
    x"365a6c36", x"3f417e3f", x"f702f5f7", x"cc4f83cc",
    x"345c6834", x"a5f451a5", x"e534d1e5", x"f108f9f1",
    x"7193e271", x"d873abd8", x"31536231", x"153f2a15",
    x"040c0804", x"c75295c7", x"23654623", x"c35e9dc3",
    x"18283018", x"96a13796", x"050f0a05", x"9ab52f9a",
    x"07090e07", x"12362412", x"809b1b80", x"e23ddfe2",
    x"eb26cdeb", x"27694e27", x"b2cd7fb2", x"759fea75",
    x"091b1209", x"839e1d83", x"2c74582c", x"1a2e341a",
    x"1b2d361b", x"6eb2dc6e", x"5aeeb45a", x"a0fb5ba0",
    x"52f6a452", x"3b4d763b", x"d661b7d6", x"b3ce7db3",
    x"297b5229", x"e33edde3", x"2f715e2f", x"84971384",
    x"53f5a653", x"d168b9d1", x"00000000", x"ed2cc1ed",
    x"20604020", x"fc1fe3fc", x"b1c879b1", x"5bedb65b",
    x"6abed46a", x"cb468dcb", x"bed967be", x"394b7239",
    x"4ade944a", x"4cd4984c", x"58e8b058", x"cf4a85cf",
    x"d06bbbd0", x"ef2ac5ef", x"aae54faa", x"fb16edfb",
    x"43c58643", x"4dd79a4d", x"33556633", x"85941185",
    x"45cf8a45", x"f910e9f9", x"02060402", x"7f81fe7f",
    x"50f0a050", x"3c44783c", x"9fba259f", x"a8e34ba8",
    x"51f3a251", x"a3fe5da3", x"40c08040", x"8f8a058f",
    x"92ad3f92", x"9dbc219d", x"38487038", x"f504f1f5",
    x"bcdf63bc", x"b6c177b6", x"da75afda", x"21634221",
    x"10302010", x"ff1ae5ff", x"f30efdf3", x"d26dbfd2",
    x"cd4c81cd", x"0c14180c", x"13352613", x"ec2fc3ec",
    x"5fe1be5f", x"97a23597", x"44cc8844", x"17392e17",
    x"c45793c4", x"a7f255a7", x"7e82fc7e", x"3d477a3d",
    x"64acc864", x"5de7ba5d", x"192b3219", x"7395e673",
    x"60a0c060", x"81981981", x"4fd19e4f", x"dc7fa3dc",
    x"22664422", x"2a7e542a", x"90ab3b90", x"88830b88",
    x"46ca8c46", x"ee29c7ee", x"b8d36bb8", x"143c2814",
    x"de79a7de", x"5ee2bc5e", x"0b1d160b", x"db76addb",
    x"e03bdbe0", x"32566432", x"3a4e743a", x"0a1e140a",
    x"49db9249", x"060a0c06", x"246c4824", x"5ce4b85c",
    x"c25d9fc2", x"d36ebdd3", x"acef43ac", x"62a6c462",
    x"91a83991", x"95a43195", x"e437d3e4", x"798bf279",
    x"e732d5e7", x"c8438bc8", x"37596e37", x"6db7da6d",
    x"8d8c018d", x"d564b1d5", x"4ed29c4e", x"a9e049a9",
    x"6cb4d86c", x"56faac56", x"f407f3f4", x"ea25cfea",
    x"65afca65", x"7a8ef47a", x"aee947ae", x"08181008",
    x"bad56fba", x"7888f078", x"256f4a25", x"2e725c2e",
    x"1c24381c", x"a6f157a6", x"b4c773b4", x"c65197c6",
    x"e823cbe8", x"dd7ca1dd", x"749ce874", x"1f213e1f",
    x"4bdd964b", x"bddc61bd", x"8b860d8b", x"8a850f8a",
    x"7090e070", x"3e427c3e", x"b5c471b5", x"66aacc66",
    x"48d89048", x"03050603", x"f601f7f6", x"0e121c0e",
    x"61a3c261", x"355f6a35", x"57f9ae57", x"b9d069b9",
    x"86911786", x"c15899c1", x"1d273a1d", x"9eb9279e",
    x"e138d9e1", x"f813ebf8", x"98b32b98", x"11332211",
    x"69bbd269", x"d970a9d9", x"8e89078e", x"94a73394",
    x"9bb62d9b", x"1e223c1e", x"87921587", x"e920c9e9",
    x"ce4987ce", x"55ffaa55", x"28785028", x"df7aa5df",
    x"8c8f038c", x"a1f859a1", x"89800989", x"0d171a0d",
    x"bfda65bf", x"e631d7e6", x"42c68442", x"68b8d068",
    x"41c38241", x"99b02999", x"2d775a2d", x"0f111e0f",
    x"b0cb7bb0", x"54fca854", x"bbd66dbb", x"163a2c16"
  );
  constant Te3 : tbox32_t := (
    x"6363a5c6", x"7c7c84f8", x"777799ee", x"7b7b8df6",
    x"f2f20dff", x"6b6bbdd6", x"6f6fb1de", x"c5c55491",
    x"30305060", x"01010302", x"6767a9ce", x"2b2b7d56",
    x"fefe19e7", x"d7d762b5", x"ababe64d", x"76769aec",
    x"caca458f", x"82829d1f", x"c9c94089", x"7d7d87fa",
    x"fafa15ef", x"5959ebb2", x"4747c98e", x"f0f00bfb",
    x"adadec41", x"d4d467b3", x"a2a2fd5f", x"afafea45",
    x"9c9cbf23", x"a4a4f753", x"727296e4", x"c0c05b9b",
    x"b7b7c275", x"fdfd1ce1", x"9393ae3d", x"26266a4c",
    x"36365a6c", x"3f3f417e", x"f7f702f5", x"cccc4f83",
    x"34345c68", x"a5a5f451", x"e5e534d1", x"f1f108f9",
    x"717193e2", x"d8d873ab", x"31315362", x"15153f2a",
    x"04040c08", x"c7c75295", x"23236546", x"c3c35e9d",
    x"18182830", x"9696a137", x"05050f0a", x"9a9ab52f",
    x"0707090e", x"12123624", x"80809b1b", x"e2e23ddf",
    x"ebeb26cd", x"2727694e", x"b2b2cd7f", x"75759fea",
    x"09091b12", x"83839e1d", x"2c2c7458", x"1a1a2e34",
    x"1b1b2d36", x"6e6eb2dc", x"5a5aeeb4", x"a0a0fb5b",
    x"5252f6a4", x"3b3b4d76", x"d6d661b7", x"b3b3ce7d",
    x"29297b52", x"e3e33edd", x"2f2f715e", x"84849713",
    x"5353f5a6", x"d1d168b9", x"00000000", x"eded2cc1",
    x"20206040", x"fcfc1fe3", x"b1b1c879", x"5b5bedb6",
    x"6a6abed4", x"cbcb468d", x"bebed967", x"39394b72",
    x"4a4ade94", x"4c4cd498", x"5858e8b0", x"cfcf4a85",
    x"d0d06bbb", x"efef2ac5", x"aaaae54f", x"fbfb16ed",
    x"4343c586", x"4d4dd79a", x"33335566", x"85859411",
    x"4545cf8a", x"f9f910e9", x"02020604", x"7f7f81fe",
    x"5050f0a0", x"3c3c4478", x"9f9fba25", x"a8a8e34b",
    x"5151f3a2", x"a3a3fe5d", x"4040c080", x"8f8f8a05",
    x"9292ad3f", x"9d9dbc21", x"38384870", x"f5f504f1",
    x"bcbcdf63", x"b6b6c177", x"dada75af", x"21216342",
    x"10103020", x"ffff1ae5", x"f3f30efd", x"d2d26dbf",
    x"cdcd4c81", x"0c0c1418", x"13133526", x"ecec2fc3",
    x"5f5fe1be", x"9797a235", x"4444cc88", x"1717392e",
    x"c4c45793", x"a7a7f255", x"7e7e82fc", x"3d3d477a",
    x"6464acc8", x"5d5de7ba", x"19192b32", x"737395e6",
    x"6060a0c0", x"81819819", x"4f4fd19e", x"dcdc7fa3",
    x"22226644", x"2a2a7e54", x"9090ab3b", x"8888830b",
    x"4646ca8c", x"eeee29c7", x"b8b8d36b", x"14143c28",
    x"dede79a7", x"5e5ee2bc", x"0b0b1d16", x"dbdb76ad",
    x"e0e03bdb", x"32325664", x"3a3a4e74", x"0a0a1e14",
    x"4949db92", x"06060a0c", x"24246c48", x"5c5ce4b8",
    x"c2c25d9f", x"d3d36ebd", x"acacef43", x"6262a6c4",
    x"9191a839", x"9595a431", x"e4e437d3", x"79798bf2",
    x"e7e732d5", x"c8c8438b", x"3737596e", x"6d6db7da",
    x"8d8d8c01", x"d5d564b1", x"4e4ed29c", x"a9a9e049",
    x"6c6cb4d8", x"5656faac", x"f4f407f3", x"eaea25cf",
    x"6565afca", x"7a7a8ef4", x"aeaee947", x"08081810",
    x"babad56f", x"787888f0", x"25256f4a", x"2e2e725c",
    x"1c1c2438", x"a6a6f157", x"b4b4c773", x"c6c65197",
    x"e8e823cb", x"dddd7ca1", x"74749ce8", x"1f1f213e",
    x"4b4bdd96", x"bdbddc61", x"8b8b860d", x"8a8a850f",
    x"707090e0", x"3e3e427c", x"b5b5c471", x"6666aacc",
    x"4848d890", x"03030506", x"f6f601f7", x"0e0e121c",
    x"6161a3c2", x"35355f6a", x"5757f9ae", x"b9b9d069",
    x"86869117", x"c1c15899", x"1d1d273a", x"9e9eb927",
    x"e1e138d9", x"f8f813eb", x"9898b32b", x"11113322",
    x"6969bbd2", x"d9d970a9", x"8e8e8907", x"9494a733",
    x"9b9bb62d", x"1e1e223c", x"87879215", x"e9e920c9",
    x"cece4987", x"5555ffaa", x"28287850", x"dfdf7aa5",
    x"8c8c8f03", x"a1a1f859", x"89898009", x"0d0d171a",
    x"bfbfda65", x"e6e631d7", x"4242c684", x"6868b8d0",
    x"4141c382", x"9999b029", x"2d2d775a", x"0f0f111e",
    x"b0b0cb7b", x"5454fca8", x"bbbbd66d", x"16163a2c"
  );
  constant Te4 : tbox8_t := (
    x"63",x"7c",x"77",x"7b",x"f2",x"6b",x"6f",x"c5",x"30",x"01",x"67",x"2b",x"fe",x"d7",x"ab",x"76",
    x"ca",x"82",x"c9",x"7d",x"fa",x"59",x"47",x"f0",x"ad",x"d4",x"a2",x"af",x"9c",x"a4",x"72",x"c0",
    x"b7",x"fd",x"93",x"26",x"36",x"3f",x"f7",x"cc",x"34",x"a5",x"e5",x"f1",x"71",x"d8",x"31",x"15",
    x"04",x"c7",x"23",x"c3",x"18",x"96",x"05",x"9a",x"07",x"12",x"80",x"e2",x"eb",x"27",x"b2",x"75",
    x"09",x"83",x"2c",x"1a",x"1b",x"6e",x"5a",x"a0",x"52",x"3b",x"d6",x"b3",x"29",x"e3",x"2f",x"84",
    x"53",x"d1",x"00",x"ed",x"20",x"fc",x"b1",x"5b",x"6a",x"cb",x"be",x"39",x"4a",x"4c",x"58",x"cf",
    x"d0",x"ef",x"aa",x"fb",x"43",x"4d",x"33",x"85",x"45",x"f9",x"02",x"7f",x"50",x"3c",x"9f",x"a8",
    x"51",x"a3",x"40",x"8f",x"92",x"9d",x"38",x"f5",x"bc",x"b6",x"da",x"21",x"10",x"ff",x"f3",x"d2",
    x"cd",x"0c",x"13",x"ec",x"5f",x"97",x"44",x"17",x"c4",x"a7",x"7e",x"3d",x"64",x"5d",x"19",x"73",
    x"60",x"81",x"4f",x"dc",x"22",x"2a",x"90",x"88",x"46",x"ee",x"b8",x"14",x"de",x"5e",x"0b",x"db",
    x"e0",x"32",x"3a",x"0a",x"49",x"06",x"24",x"5c",x"c2",x"d3",x"ac",x"62",x"91",x"95",x"e4",x"79",
    x"e7",x"c8",x"37",x"6d",x"8d",x"d5",x"4e",x"a9",x"6c",x"56",x"f4",x"ea",x"65",x"7a",x"ae",x"08",
    x"ba",x"78",x"25",x"2e",x"1c",x"a6",x"b4",x"c6",x"e8",x"dd",x"74",x"1f",x"4b",x"bd",x"8b",x"8a",
    x"70",x"3e",x"b5",x"66",x"48",x"03",x"f6",x"0e",x"61",x"35",x"57",x"b9",x"86",x"c1",x"1d",x"9e",
    x"e1",x"f8",x"98",x"11",x"69",x"d9",x"8e",x"94",x"9b",x"1e",x"87",x"e9",x"ce",x"55",x"28",x"df",
    x"8c",x"a1",x"89",x"0d",x"bf",x"e6",x"42",x"68",x"41",x"99",x"2d",x"0f",x"b0",x"54",x"bb",x"16"
  );

  -- Inverse S-box Td4
  constant Td4 : tbox8_t := (
    x"52",x"09",x"6a",x"d5",x"30",x"36",x"a5",x"38",x"bf",x"40",x"a3",x"9e",x"81",x"f3",x"d7",x"fb",
    x"7c",x"e3",x"39",x"82",x"9b",x"2f",x"ff",x"87",x"34",x"8e",x"43",x"44",x"c4",x"de",x"e9",x"cb",
    x"54",x"7b",x"94",x"32",x"a6",x"c2",x"23",x"3d",x"ee",x"4c",x"95",x"0b",x"42",x"fa",x"c3",x"4e",
    x"08",x"2e",x"a1",x"66",x"28",x"d9",x"24",x"b2",x"76",x"5b",x"a2",x"49",x"6d",x"8b",x"d1",x"25",
    x"72",x"f8",x"f6",x"64",x"86",x"68",x"98",x"16",x"d4",x"a4",x"5c",x"cc",x"5d",x"65",x"b6",x"92",
    x"6c",x"70",x"48",x"50",x"fd",x"ed",x"b9",x"da",x"5e",x"15",x"46",x"57",x"a7",x"8d",x"9d",x"84",
    x"90",x"d8",x"ab",x"00",x"8c",x"bc",x"d3",x"0a",x"f7",x"e4",x"58",x"05",x"b8",x"b3",x"45",x"06",
    x"d0",x"2c",x"1e",x"8f",x"ca",x"3f",x"0f",x"02",x"c1",x"af",x"bd",x"03",x"01",x"13",x"8a",x"6b",
    x"3a",x"91",x"11",x"41",x"4f",x"67",x"dc",x"ea",x"97",x"f2",x"cf",x"ce",x"f0",x"b4",x"e6",x"73",
    x"96",x"ac",x"74",x"22",x"e7",x"ad",x"35",x"85",x"e2",x"f9",x"37",x"e8",x"1c",x"75",x"df",x"6e",
    x"47",x"f1",x"1a",x"71",x"1d",x"29",x"c5",x"89",x"6f",x"b7",x"62",x"0e",x"aa",x"18",x"be",x"1b",
    x"fc",x"56",x"3e",x"4b",x"c6",x"d2",x"79",x"20",x"9a",x"db",x"c0",x"fe",x"78",x"cd",x"5a",x"f4",
    x"1f",x"dd",x"a8",x"33",x"88",x"07",x"c7",x"31",x"b1",x"12",x"10",x"59",x"27",x"80",x"ec",x"5f",
    x"60",x"51",x"7f",x"a9",x"19",x"b5",x"4a",x"0d",x"2d",x"e5",x"7a",x"9f",x"93",x"c9",x"9c",x"ef",
    x"a0",x"e0",x"3b",x"4d",x"ae",x"2a",x"f5",x"b0",x"c8",x"eb",x"bb",x"3c",x"83",x"53",x"99",x"61",
    x"17",x"2b",x"04",x"7e",x"ba",x"77",x"d6",x"26",x"e1",x"69",x"14",x"63",x"55",x"21",x"0c",x"7d"
  );
  -- TODO: populate Td0..Td3 if decryption core needs table-based rounds
  constant Td0 : tbox32_t := (others => (others => '0'));
  constant Td1 : tbox32_t := (others => (others => '0'));
  constant Td2 : tbox32_t := (others => (others => '0'));
  constant Td3 : tbox32_t := (others => (others => '0'));

end package body;

